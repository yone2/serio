`timescale 1ns/1ps

module case_rom(romaddr, t_cmd, t_addr, t_data);
input  [7:0] romaddr;
output [1:0] t_cmd;
output [7:0] t_addr;
output [7:0] t_data;

assign {t_cmd, t_addr, t_data} = rom_table(romaddr);

function [17:0] rom_table;
	input addr;
	case (addr)
	8'h00   : rom_table = 18'h1_01_40;
	8'h01   : rom_table = 18'h1_02_60;
	8'h02   : rom_table = 18'h1_03_0a;
	8'h03   : rom_table = 18'h1_0c_00;
	8'h04   : rom_table = 18'h1_0e_61;
	8'h05   : rom_table = 18'h1_0f_4b;
	8'h06   : rom_table = 18'h1_15_00;
	8'h07   : rom_table = 18'h1_16_02;
	8'h08   : rom_table = 18'h1_17_13;
	8'h09   : rom_table = 18'h1_18_01;
	8'h0a   : rom_table = 18'h1_19_02;
	8'h0b   : rom_table = 18'h1_1a_7a;
	8'h0c   : rom_table = 18'h1_1e_07;
	8'h0d   : rom_table = 18'h1_21_02;
	8'h0e   : rom_table = 18'h1_22_91;
	8'h0f   : rom_table = 18'h1_29_07;
	8'h10   : rom_table = 18'h1_32_b6;
	8'h11   : rom_table = 18'h1_33_0b;
	8'h12   : rom_table = 18'h1_34_11;
	8'h13   : rom_table = 18'h1_35_0b;
	8'h14   : rom_table = 18'h1_37_1d;
	8'h15   : rom_table = 18'h1_38_71;
	8'h16   : rom_table = 18'h1_39_2a;
	8'h17   : rom_table = 18'h1_3b_12;
	8'h18   : rom_table = 18'h1_3c_78;
	8'h19   : rom_table = 18'h1_3d_c3;
	8'h1a   : rom_table = 18'h1_3e_00;
	8'h1b   : rom_table = 18'h1_3f_00;
	8'h1c   : rom_table = 18'h1_41_08; // ?
	8'h1d   : rom_table = 18'h1_41_38;
	8'h1e   : rom_table = 18'h1_43_0a;
	8'h1f   : rom_table = 18'h1_44_f0;
	8'h20   : rom_table = 18'h1_45_34;
	8'h21   : rom_table = 18'h1_46_58;
	8'h22   : rom_table = 18'h1_47_28;
	8'h23   : rom_table = 18'h1_48_3a;
	8'h24   : rom_table = 18'h1_4b_09;
	8'h25   : rom_table = 18'h1_4c_00;
	8'h26   : rom_table = 18'h1_4d_40;
	8'h27   : rom_table = 18'h1_4e_20;
	8'h28   : rom_table = 18'h1_4f_80;
	8'h29   : rom_table = 18'h1_50_80;
	8'h2a   : rom_table = 18'h1_51_00;
	8'h2b   : rom_table = 18'h1_52_22;
	8'h2c   : rom_table = 18'h1_53_5e;
	8'h2d   : rom_table = 18'h1_54_80;
	8'h2e   : rom_table = 18'h1_56_40;
	8'h2f   : rom_table = 18'h1_58_9e;
	8'h30   : rom_table = 18'h1_59_88;
	8'h31   : rom_table = 18'h1_5a_88;
	8'h32   : rom_table = 18'h1_5b_44;
	8'h33   : rom_table = 18'h1_5c_67;
	8'h34   : rom_table = 18'h1_5d_49;
	8'h35   : rom_table = 18'h1_5e_0e;
	8'h36   : rom_table = 18'h1_69_00;
	8'h37   : rom_table = 18'h1_6a_40;
	8'h38   : rom_table = 18'h1_6b_0a;
	8'h39   : rom_table = 18'h1_6c_0a;
	8'h3a   : rom_table = 18'h1_6d_55;
	8'h3b   : rom_table = 18'h1_6e_11;
	8'h3c   : rom_table = 18'h1_6f_9f;
	8'h3d   : rom_table = 18'h1_70_3a;
	8'h3e   : rom_table = 18'h1_71_35;
	8'h3f   : rom_table = 18'h1_72_11;
	8'h40   : rom_table = 18'h1_73_f0;
	8'h41   : rom_table = 18'h1_74_10;
	8'h42   : rom_table = 18'h1_75_05;
	8'h43   : rom_table = 18'h1_76_e1;
	8'h44   : rom_table = 18'h1_77_01;
	8'h45   : rom_table = 18'h1_78_04;
	8'h46   : rom_table = 18'h1_79_01;
	8'h47   : rom_table = 18'h1_8d_4f;
	8'h48   : rom_table = 18'h1_8e_00;
	8'h49   : rom_table = 18'h1_8f_00;
	8'h4a   : rom_table = 18'h1_90_00;
	8'h4b   : rom_table = 18'h1_91_00;
	8'h4c   : rom_table = 18'h1_96_00;
	8'h4d   : rom_table = 18'h1_96_00;
	8'h4e   : rom_table = 18'h1_97_30;
	8'h4f   : rom_table = 18'h1_98_20;
	8'h50   : rom_table = 18'h1_99_30;
	8'h51   : rom_table = 18'h1_9a_00;
	8'h52   : rom_table = 18'h1_9a_84;
	8'h53   : rom_table = 18'h1_9b_29;
	8'h54   : rom_table = 18'h1_9c_03;
	8'h55   : rom_table = 18'h1_9d_4c;
	8'h56   : rom_table = 18'h1_9e_3f;
	8'h57   : rom_table = 18'h1_a2_02;
	8'h58   : rom_table = 18'h1_a4_88;
	8'h59   : rom_table = 18'h1_b0_84;
	8'h5a   : rom_table = 18'h1_b1_0c;
	8'h5b   : rom_table = 18'h1_b2_0e;
	8'h5c   : rom_table = 18'h1_b3_82;
	8'h5d   : rom_table = 18'h1_b8_0a;
	8'h5e   : rom_table = 18'h1_c8_f0;
	8'h5f   : rom_table = 18'h1_c9_60;
	default : rom_table = 18'h1_00_00;
	endcase
endfunction

endmodule
